library ieee;
use ieee.std_logic_1164.all;
use work.std_arith.all;

use work.paquete.all;

entity tabletBottlingSystem is

end tabletBottlingSystem;

architecture funcional of tabletBottlingSystem is

end funcional;